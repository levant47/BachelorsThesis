package program is
    constant code : work.types.T_MEMORY := (
        b"00000001",
        b"00000000",
        b"00001100",
        b"00000001",
        b"00000001",
        b"00000100",
        b"00000111",
        b"00001010",
        b"00001011",
        b"00010100",
        b"00000001",
        b"00000000",
        b"00000001",
        b"00000001",
        b"00001101",
        b"00000010",
        b"00000001",
        b"00000000",
        b"00001011",
        b"00011100",
        b"00000001",
        b"00000000",
        b"00000001",
        b"00000000",
        b"00001101",
        b"00000010",
        b"00000001",
        b"00000001",
        b"00000001",
        b"01100100",
        b"00001100",
        b"00000001",
        b"00000000",
        b"00000100",
        b"00000111",
        b"01000101",
        b"00000001",
        b"01100100",
        b"00001100",
        b"00000001",
        b"00000000",
        b"00000100",
        b"00000111",
        b"00111111",
        b"00000001",
        b"01100100",
        b"00001100",
        b"00000001",
        b"00000000",
        b"00000100",
        b"00000111",
        b"00111001",
        b"00000001",
        b"11111111",
        b"00000011",
        b"00001011",
        b"00101110",
        b"00000010",
        b"00000001",
        b"11111111",
        b"00000011",
        b"00001011",
        b"00100110",
        b"00000010",
        b"00000001",
        b"11111111",
        b"00000011",
        b"00001011",
        b"00011110",
        b"00000010",
        b"00001011",
        b"00000010"
    );
end program;
