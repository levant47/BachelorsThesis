library IEEE;
use IEEE.std_logic_1164.all;
package program is
    constant code : work.types.T_MEMORY := (
        b"00000001",
        b"00000001",
        b"00010000",
        b"00000001",
        b"00000000",
        b"00010001",
        b"00001100",
        b"00010000",
        b"00001101",
        b"00000001",
        b"00110010",
        b"00000001",
        b"11011100",
        b"00000001",
        b"11010101",
        b"00000001",
        b"01001110",
        b"00000001",
        b"00010101",
        b"00010000",
        b"00001011",
        b"00010001",
        b"00000001",
        b"01101110",
        b"00000001",
        b"00011100",
        b"00010000",
        b"00001011",
        b"00010000",
        b"00000001",
        b"00000011",
        b"00001011",
        b"00001100",
        b"00000001",
        b"00000000",
        b"00000100",
        b"00000001",
        b"00101101",
        b"00000111",
        b"00000001",
        b"11111111",
        b"00000011",
        b"00000001",
        b"00100000",
        b"00001011",
        b"00000010",
        b"00010001",
        b"00001011",
        b"00000001",
        b"00100000",
        b"00000001",
        b"00110110",
        b"00010000",
        b"00001011",
        b"00001100",
        b"00000001",
        b"00000000",
        b"00000100",
        b"00000001",
        b"01001011",
        b"00000111",
        b"00000001",
        b"11111111",
        b"00000001",
        b"00100000",
        b"00000001",
        b"01000101",
        b"00010000",
        b"00001011",
        b"00000001",
        b"11111111",
        b"00000011",
        b"00000001",
        b"00110110",
        b"00001011",
        b"00000010",
        b"00010001",
        b"00001011",
        b"00000001",
        b"00110000",
        b"00000001",
        b"01010100",
        b"00010000",
        b"00001011",
        b"00001100",
        b"00000001",
        b"00000000",
        b"00000100",
        b"00000001",
        b"01101011",
        b"00000111",
        b"00000001",
        b"11111111",
        b"00000001",
        b"11111111",
        b"00000001",
        b"00110000",
        b"00000001",
        b"01100101",
        b"00010000",
        b"00001011",
        b"00000001",
        b"11111111",
        b"00000011",
        b"00000001",
        b"01010100",
        b"00001011",
        b"00000010",
        b"00010001",
        b"00001011",
        b"00000001",
        b"00000000",
        b"00000100",
        b"00000001",
        b"01111000",
        b"00000111",
        b"00000001",
        b"00000000",
        b"00010001",
        b"00001011",
        b"00000001",
        b"00000001",
        b"00010001",
        b"00001011"
    );
end program;
