library IEEE;
use IEEE.std_logic_1164.all;
package program is
    constant code : work.types.T_MEMORY := (
        b"00001110",
        b"00001110",
        b"00001110",
        b"00000001",
        b"00000011",
        b"00001011"
    );
end program;
