library IEEE;
use IEEE.std_logic_1164.all;
package program is
    constant code : work.types.T_MEMORY := (
        b"00000001",
        b"00001010",
        b"00001100",
        b"00000001",
        b"00000000",
        b"00000100",
        b"00000001",
        b"00001111",
        b"00000111",
        b"00000001",
        b"11111111",
        b"00000011",
        b"00000001",
        b"00000010",
        b"00001011",
        b"00000010",
        b"00000001",
        b"00010000",
        b"00001011"
    );
end program;
